image/svg+xml;charset=UTF-8,%3csvg width='4' height='4' viewBox='0 0 4 4' fill='none' xmlns='http://www.w3.org/2000/svg'%3e%3ccircle cx='2' cy='2' r='2' fill='%23FF532E'/%3e%3c/svg%3e